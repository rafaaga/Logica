-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri May 27 18:31:18 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY matrizLeds IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        R0 : OUT STD_LOGIC;
        R1 : OUT STD_LOGIC;
        R2 : OUT STD_LOGIC;
        R3 : OUT STD_LOGIC;
        R4 : OUT STD_LOGIC;
        R5 : OUT STD_LOGIC;
        R6 : OUT STD_LOGIC;
        R7 : OUT STD_LOGIC
    );
END matrizLeds;

ARCHITECTURE BEHAVIOR OF matrizLeds IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6,state7,state8);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            R0 <= '0';
            R1 <= '0';
            R2 <= '0';
            R3 <= '0';
            R4 <= '0';
            R5 <= '0';
            R6 <= '0';
            R7 <= '0';
        ELSE
            R0 <= '0';
            R1 <= '0';
            R2 <= '0';
            R3 <= '0';
            R4 <= '0';
            R5 <= '0';
            R6 <= '0';
            R7 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    reg_fstate <= state2;

                    R0 <= '1';

                    R7 <= '0';

                    R6 <= '0';

                    R5 <= '0';

                    R4 <= '0';

                    R3 <= '0';

                    R2 <= '0';

                    R1 <= '0';
                WHEN state2 =>
                    reg_fstate <= state3;

                    R0 <= '0';

                    R7 <= '0';

                    R6 <= '0';

                    R5 <= '0';

                    R4 <= '0';

                    R3 <= '0';

                    R2 <= '0';

                    R1 <= '1';
                WHEN state3 =>
                    reg_fstate <= state4;

                    R0 <= '0';

                    R7 <= '0';

                    R6 <= '0';

                    R5 <= '0';

                    R4 <= '0';

                    R3 <= '0';

                    R2 <= '1';

                    R1 <= '0';
                WHEN state4 =>
                    reg_fstate <= state5;

                    R0 <= '0';

                    R7 <= '0';

                    R6 <= '0';

                    R5 <= '0';

                    R4 <= '0';

                    R3 <= '1';

                    R2 <= '0';

                    R1 <= '0';
                WHEN state5 =>
                    reg_fstate <= state6;

                    R0 <= '0';

                    R7 <= '0';

                    R6 <= '0';

                    R5 <= '0';

                    R4 <= '1';

                    R3 <= '0';

                    R2 <= '0';

                    R1 <= '0';
                WHEN state6 =>
                    reg_fstate <= state7;

                    R0 <= '0';

                    R7 <= '0';

                    R6 <= '0';

                    R5 <= '1';

                    R4 <= '0';

                    R3 <= '0';

                    R2 <= '0';

                    R1 <= '0';
                WHEN state7 =>
                    reg_fstate <= state8;

                    R0 <= '0';

                    R7 <= '0';

                    R6 <= '1';

                    R5 <= '0';

                    R4 <= '0';

                    R3 <= '0';

                    R2 <= '0';

                    R1 <= '0';
                WHEN state8 =>
                    reg_fstate <= state1;

                    R0 <= '0';

                    R7 <= '1';

                    R6 <= '0';

                    R5 <= '0';

                    R4 <= '0';

                    R3 <= '0';

                    R2 <= '0';

                    R1 <= '0';
                WHEN OTHERS => 
                    R0 <= 'X';
                    R1 <= 'X';
                    R2 <= 'X';
                    R3 <= 'X';
                    R4 <= 'X';
                    R5 <= 'X';
                    R6 <= 'X';
                    R7 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
